--
-- CycleController.vhd
--
-- Finite-state machine to control the wash cycles of a washing machine.
--
-- ELEE 204 Design Project
--   Kaleb Dekker, JD Elsey, David Fritts, Domenic Rodriguez
--
-- April 12, 2016 
--

-- Import required libraries
library IEEE;
use IEEE.std_logic_1164.all;

entity CycleController is

end;

architecture CycleController_arch of CycleController is
begin

end CycleController_arch;
