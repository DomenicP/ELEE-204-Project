--
-- PaymentController.vhd
--
-- Finite-state machine to control payments for a washing machine.
--
-- ELEE 204 Design Project
--   Kaleb Dekker, JD Elsey, David Fritts, Domenic Rodriguez
--
-- April 12, 2016 
--

-- Import required libraries
library IEEE;
use IEEE.std_logic_1164.all;

entity PaymentController is

end PaymentController;

architecture PaymentController_arch of PaymentController is
begin

end PaymentController_arch;
